module MAR(input clk, input ld, wr, rst, input [31:0] PC, output [31:0] address);

endmodule 

module memory(input [31:0] address, output [31:0] data)

endmodule

module MDR(input clk, input ld, wr, rst, input [31:0] data_in, output [31:0] data_out);

endmodule 