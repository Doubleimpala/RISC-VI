module cpu_core(input clk, input rst);


endmodule